module rc4_tb();
    reg 
endmodule 