module rc4_inst();

endmodule